** Profile: "SCHEMATIC1-lab3r"  [ D:\academic glasgow\junior second\ccd\labfile\lab3-pspicefiles\schematic1\lab3r.sim ] 

** Creating circuit file "lab3r.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
.INC "D:\academic glasgow\junior second\ccd\labfile\lab3-pspicefiles\schematic1\lab3r\lab3r_profile.inc" 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\Amberisy\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 50ms 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
